module testBench()

endmodule